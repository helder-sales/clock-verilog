//Debouncer
module debouncer(input in, clk, output reg out);

reg op1, op2, op3;

/*------------------------------------------------------------------------------------*/

always @(posedge clk)
	begin
	
		op1 = in;

		op2 = op1;

		op3 = op2;	

		out <= op1 & op2 & op3;
	
	end
	
endmodule 

/*------------------------------------------------------------------------------------
  ------------------------------------------------------------------------------------*/